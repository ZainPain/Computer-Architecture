library verilog;
use verilog.vl_types.all;
entity truncator_sv_unit is
end truncator_sv_unit;
