library verilog;
use verilog.vl_types.all;
entity cache_arbiter_sv_unit is
end cache_arbiter_sv_unit;
