library verilog;
use verilog.vl_types.all;
entity or_sv_unit is
end or_sv_unit;
