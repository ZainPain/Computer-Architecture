library verilog;
use verilog.vl_types.all;
entity IF_ID_reg_sv_unit is
end IF_ID_reg_sv_unit;
