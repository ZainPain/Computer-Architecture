library verilog;
use verilog.vl_types.all;
entity Hazard20Detection_sv_unit is
end Hazard20Detection_sv_unit;
