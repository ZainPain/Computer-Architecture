library verilog;
use verilog.vl_types.all;
entity extract_cache_components_sv_unit is
end extract_cache_components_sv_unit;
