library verilog;
use verilog.vl_types.all;
entity Address_checker_sv_unit is
end Address_checker_sv_unit;
