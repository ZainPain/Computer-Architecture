library verilog;
use verilog.vl_types.all;
entity NOPS_sv_unit is
end NOPS_sv_unit;
