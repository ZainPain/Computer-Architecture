library verilog;
use verilog.vl_types.all;
entity adj_imm_sv_unit is
end adj_imm_sv_unit;
