library verilog;
use verilog.vl_types.all;
entity ID_EX_reg_sv_unit is
end ID_EX_reg_sv_unit;
