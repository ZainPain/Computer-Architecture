library verilog;
use verilog.vl_types.all;
entity memory_caches_sv_unit is
end memory_caches_sv_unit;
