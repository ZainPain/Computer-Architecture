library verilog;
use verilog.vl_types.all;
entity LRU_register_sv_unit is
end LRU_register_sv_unit;
