library verilog;
use verilog.vl_types.all;
entity \__and___sv_unit\ is
end \__and___sv_unit\;
