library verilog;
use verilog.vl_types.all;
entity writeback_forward_sv_unit is
end writeback_forward_sv_unit;
