import lc3b_types::*;
module cache_datapath
(
)

endmodule cache_datapath