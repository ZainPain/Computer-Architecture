library verilog;
use verilog.vl_types.all;
entity MEM_WB_reg_sv_unit is
end MEM_WB_reg_sv_unit;
