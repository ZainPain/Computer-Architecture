library verilog;
use verilog.vl_types.all;
entity mask_sv_unit is
end mask_sv_unit;
