library verilog;
use verilog.vl_types.all;
entity \_8by1mux_sv_unit\ is
end \_8by1mux_sv_unit\;
