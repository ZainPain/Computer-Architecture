library verilog;
use verilog.vl_types.all;
entity Memory_mapped_IO_sv_unit is
end Memory_mapped_IO_sv_unit;
