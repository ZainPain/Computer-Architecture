library verilog;
use verilog.vl_types.all;
entity staller_sv_unit is
end staller_sv_unit;
