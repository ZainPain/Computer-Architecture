library verilog;
use verilog.vl_types.all;
entity write_to_dataArray_sv_unit is
end write_to_dataArray_sv_unit;
