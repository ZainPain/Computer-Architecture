library verilog;
use verilog.vl_types.all;
entity Forwarding_sv_unit is
end Forwarding_sv_unit;
